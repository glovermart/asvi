// NOTE: Line 13.

interface I;

  logic x;

endinterface


module top; 
  
   struct
    { I u_I; // Parenthesis omitted.
    } st_Ifc;

endmodule
