module tb;
 top u_DUT();
 initial begin
  $info("Testing Simulation of Initial Testcases");
  $finish;
 end
endmodule
