// Assignment via `always_latch` to scalar members of an SVI port.
// Array of SVIs

// Using modports, output 'y' from module M1 is an input to module M2.

/* Modules M1 and M2 now with en and arst pins connected directly to 
 top module pins.*/

/* Removed nets not used in modport to avoid inferred connection to 
 to the input or output of other module (M1 or M2).*/


`define V 8

interface I;
  timeunit 1ns;
  timeprecision 1ps;
  
  logic y;

  modport P1
    ( 
     output y
    );

  modport P2
    ( input y
    );

endinterface

module M1
  ( I.P1 p1[`V-1:0]
  , output logic [`V-1:0]o_a
  , input logic en
  , input logic i_arst
  );
  timeunit 1ns;
  timeprecision 1ps;
  
  for(genvar i =0; i< `V;i++) begin
    always_latch begin
      if (!i_arst)
        p1[i].y <= 1'b0;
      else if (en)
        p1[i].y <= 1'b1;
    end
  assign o_a[i] = p1[i].y;
  end

endmodule

/* A different enable signal may be used in M2 to make en
 independent */ 
 
module M2
  ( I.P2 p2[`V-1:0]
  , output logic [`V-1:0]o_b
  , input logic en
  );
  timeunit 1ns;
  timeprecision 1ps;

  for(genvar i =0; i< `V;i++) begin
    always_latch begin
     if (en)
       o_b[i] <= p2[i].y;
    end
  end

endmodule



module top
  ( input logic en
  , input logic i_clk
  , input logic i_arst
  , output logic [`V-1:0]o_a 
  , output logic [`V-1:0]o_b
  );

  timeunit 1ns;
  timeprecision 1ps;
  
  I u_I [`V-1:0] ();

  M1 u_M1
    ( .p1(u_I)
    , .o_a(o_a)
    , .en
    , .i_arst 
    );

  M2 u_M2
    ( .p2(u_I)
    , .o_b(o_b)
    , .en
    );

endmodule
